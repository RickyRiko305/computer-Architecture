library verilog;
use verilog.vl_types.all;
entity Block3_vlg_vec_tst is
end Block3_vlg_vec_tst;
