library verilog;
use verilog.vl_types.all;
entity alu_bcd_vlg_vec_tst is
end alu_bcd_vlg_vec_tst;
