library verilog;
use verilog.vl_types.all;
entity ALU_32_bit_vlg_vec_tst is
end ALU_32_bit_vlg_vec_tst;
