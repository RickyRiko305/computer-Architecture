library verilog;
use verilog.vl_types.all;
entity q1_1_vlg_vec_tst is
end q1_1_vlg_vec_tst;
