library verilog;
use verilog.vl_types.all;
entity Block4_vlg_vec_tst is
end Block4_vlg_vec_tst;
