library verilog;
use verilog.vl_types.all;
entity Block3_vlg_check_tst is
    port(
        g               : in     vl_logic;
        h               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Block3_vlg_check_tst;
