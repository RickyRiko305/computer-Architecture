library verilog;
use verilog.vl_types.all;
entity ALU32_vlg_vec_tst is
end ALU32_vlg_vec_tst;
