library verilog;
use verilog.vl_types.all;
entity bcd_7_segment_vlg_vec_tst is
end bcd_7_segment_vlg_vec_tst;
