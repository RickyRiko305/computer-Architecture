library verilog;
use verilog.vl_types.all;
entity Block3 is
    port(
        g               : out    vl_logic;
        w1              : in     vl_logic;
        w2              : in     vl_logic;
        w3              : in     vl_logic;
        w4              : in     vl_logic;
        h               : out    vl_logic
    );
end Block3;
