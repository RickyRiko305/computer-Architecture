library verilog;
use verilog.vl_types.all;
entity Lab1_1_vlg_vec_tst is
end Lab1_1_vlg_vec_tst;
