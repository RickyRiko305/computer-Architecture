library verilog;
use verilog.vl_types.all;
entity Block3_vlg_sample_tst is
    port(
        w1              : in     vl_logic;
        w2              : in     vl_logic;
        w3              : in     vl_logic;
        w4              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Block3_vlg_sample_tst;
