library verilog;
use verilog.vl_types.all;
entity q2_pc_vlg_vec_tst is
end q2_pc_vlg_vec_tst;
