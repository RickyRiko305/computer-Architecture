library verilog;
use verilog.vl_types.all;
entity verfunctions_vlg_vec_tst is
end verfunctions_vlg_vec_tst;
